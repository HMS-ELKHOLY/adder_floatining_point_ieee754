library verilog;
use verilog.vl_types.all;
entity t is
end t;
